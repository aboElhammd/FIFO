package shared_package;
	int error_count=0;
	int correct_count=0;
	bit test_finished;
endpackage : shared_package
